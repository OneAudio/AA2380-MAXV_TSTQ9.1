CONSTVAL_inst : CONSTVAL PORT MAP (
		result	 => result_sig
	);
